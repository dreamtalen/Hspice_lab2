.TITLE Adder_Top
.lib "/home/wjin/dmtalen/hspice/Hspice_lab1/PTM/models" ptm16lstp
.options acct list post
.global vdd gnd vss
.TEMP 85
.param h=4
.param vds_sup=0.1
.param SUPPLY=0.85
.param supplyB=0

.param finp=2
.param finn=1
.param length=20n
.param fint=12n
.param finh=26n

.param D=1

.param H1=1
.param H2=1
.param H3=1
.param H4=1
.param H5=1
.param H6=1
.param H7=1
.param H8=1
.param HINV=10
*********************Sub model************
*********************INV************
.SUBCKT INV A Y nfinn=2 nfinp=2
xnmos Y A GND GND lnfet l=length nfin=nfinn
xpmos Y A VDD VDD lpfet l=length nfin=nfinp
.ENDS
*********************PROP************
.SUBCKT PROP ai bi aib bib clk pi nfinn=30 nfinp=30
xnmos1 A clk GND GND lnfet l=length nfin=nfinn
xnmos2 B ai A GND lnfet l=length nfin=nfinn
xnmos3 D bib B GND lnfet l=length nfin=nfinn
xnmos4 C bi A GND lnfet l=length nfin=nfinn
xnmos5 D aib C GND lnfet l=length nfin=nfinn

xpmos1 D clk VDD VDD lpfet l=length nfin=2
xpmos2 D E VDD VDD lpfet l=length nfin=2
X1 D E INV
X2 D pi INV
.ENDS
*********************GENERATE************
.SUBCKT GENERATE A B CLK G nfinn=30 nfinp=10
xpmos1 C CLK VDD VDD lpfet l=length nfin=nfinp
xpmos2 C F VDD VDD lpfet l=length nfin=nfinp

X_INV1 C F INV

xnmos1 C A D GND lnfet l=length nfin=nfinn
xnmos2 D B E GND lnfet l=length nfin=nfinn
xnmos3 E CLK GND GND lnfet l=length nfin=nfinn

X_INV2 C G INV

.ENDS
*********************DOT_G************
.SUBCKT Dot_G Gi1 Gi2 Pi2 clk Gout nfinn=10 nfinp=30
xnmos1 A Gi1 GND GND lnfet l=length nfin=nfinn
xnmos2 B Pi2 A GND lnfet l=length nfin=nfinn
xnmos3 B Gi2 GND GND lnfet l=length nfin=nfinn

xpmos1 B clk VDD VDD lpfet l=length nfin=nfinp
xpmos2 B C VDD VDD lpfet l=length nfin=5                                                                                      
X1 B C INV
X2 B Gout INV
.ENDS
*********************DOT_P************
.SUBCKT DOT_P P1 P2 CLK P_OUT nfinn=30 nfinp=10
xpmos1 A CLK VDD VDD lpfet l=length nfin=nfinp
xpmos2 A C VDD VDD lpfet l=length nfin=nfinp

X_INV1 A C INV

xnmos1 A P1 B GND lnfet l=length nfin=nfinn
xnmos2 B P2 GND GND lnfet l=length nfin=nfinn

X_INV2 A P_OUT INV

.ENDS
*********************DOT************
.SUBCKT DOT Gi1 Pi1 Gi2 Pi2 Gout Pout CLK
XDot_G Gi1 Gi2 Pi2 clk Gout DOT_G
XDot_P Pi1 Pi2 clk Pout DOT_P
.ENDS
*********************SUM************
.SUBCKT SUM  S0 S1 C_IN CLK CLK_D SUM_OUT nfinn=30 nfinp=10
xpmos1 A CLK VDD VDD lpfet l=length nfin=40
xnmos1 A C_IN B GND lnfet l=length nfin=5
xnmos2 B CLK GND GND lnfet l=length nfin=5

xpmos2 C CLK VDD VDD lpfet l=length nfin=nfinp
xnmos3 C C_IN D GND lnfet l=length nfin=nfinn
xnmos4 D S1 E GND lnfet l=length nfin=nfinn
xnmos5 E CLK GND GND lnfet l=length nfin=nfinn

xpmos3 F CLK_D VDD VDD lpfet l=length nfin=nfinp
xpmos4 F G VDD VDD lpfet l=length nfin=2
X_INV1 F G INV
xnmos6 F A H GND lnfet l=length nfin=10
xnmos7 H S0 I GND lnfet l=length nfin=50
xnmos8 I CLK_D GND GND lnfet l=length nfin=50

xpmos5 SUM_OUT F VDD VDD lpfet l=length nfin=nfinp
xnmos9 SUM_OUT F J GND lnfet l=length nfin=nfinn
xnmos10 J C GND GND lnfet l=length nfin=nfinn
xpmos6 SUM_OUT C VDD VDD lpfet l=length nfin=nfinp

.ENDS
*********************CLK Chain For Five Level************
.SUBCKT CLKChain CLK CLKNEXT nfinn=20 nfinp=20
XCLKINV1 CLK A INV M='2'
xpmos5 B GND A VDD lpfet l=length nfin=nfinp
xnmos9 A VDD B GND lnfet l=length nfin=nfinn
XCLKINV2 B CLKNEXT INV M='2'
.ENDS

*********************CLK Delay************
.SUBCKT CLKDelay CLK CLKD nfinn=2 nfinp=2
XCLKINV1 CLK A INV M='10'
xpmos5 B GND A VDD lpfet l=length nfin=nfinp
xnmos9 A VDD B GND lnfet l=length nfin=nfinn
XCLKINV2 B CLKD INV M='10'
.ENDS
*********************TOP Circuit**********
*********************CLK Delayed Domino************
*XCLK0  CLK  CLK1  CLKChain
*XCLK1  CLK1  CLK2  CLKChain
*XCLK2  CLK2  CLK3  CLKChain
*XCLK3  CLK3  CLK4  CLKChain
*XCLK4  CLK4  CLK5  CLKChain
*XCLK5  CLK5  CLK6  CLKChain

*XCLK1D  CLK1  CLK1_D  CLKDelay
*XCLK2D  CLK2  CLK2_D  CLKDelay
*XCLK3D1  CLK  CLK_D  CLKDelay
*XCLK3D2  CLK_D1  CLK_D2  CLKDelay
*XCLK3D3  CLK_D2  CLK_D  CLKDelay
*XCLK3D4  CLK_D3  CLK_D4  CLKDelay
*XCLK3D5  CLK_D4  CLK_D5  CLKDelay
*XCLK3D6  CLK_D5  CLK_D6  CLKDelay
*XCLK3D7  CLK_D6  CLK_D  CLKDelay

*********************Inverse Signal**********
     ********************Inverse A**********
XP0Ab  A0  A0B  INV
XP1Ab  A1  A1B  INV
XP2Ab  A2  A2B  INV
XP3Ab  A3  A3B  INV
XP4Ab  A4  A4B  INV
XP5Ab  A5  A5B  INV
XP6Ab  A6  A6B  INV
XP7Ab  A7  A7B  INV
XP8Ab  A8  A8B  INV
XP9Ab  A9  A9B  INV
XP10Ab  A10  A10B  INV
XP11Ab  A11  A11B  INV
XP12Ab  A12  A12B  INV
XP13Ab  A13  A13B  INV
XP14Ab  A14  A14B  INV
XP15Ab  A15  A15B  INV
XP16Ab  A16  A16B  INV
XP17Ab  A17  A17B  INV
XP18Ab  A18  A18B  INV
XP19Ab  A19  A19B  INV
XP20Ab  A20  A20B  INV
XP21Ab  A21  A21B  INV
XP22Ab  A22  A22B  INV
XP23Ab  A23  A23B  INV
XP24Ab  A24  A24B  INV
XP25Ab  A25  A25B  INV
XP26Ab  A26  A26B  INV
XP27Ab  A27  A27B  INV
XP28Ab  A28  A28B  INV
XP29Ab  A29  A29B  INV
XP30Ab  A30  A30B  INV
XP31Ab  A31  A31B  INV
      ********************Inverse B**********
XP0Bb  B0  B0B  INV
XP1Bb  B1  B1B  INV
XP2Bb  B2  B2B  INV
XP3Bb  B3  B3B  INV
XP4Bb  B4  B4B  INV
XP5Bb  B5  B5B  INV
XP6Bb  B6  B6B  INV
XP7Bb  B7  B7B  INV
XP8Bb  B8  B8B  INV
XP9Bb  B9  B9B  INV
XP10Bb  B10  B10B  INV
XP11Bb  B11  B11B  INV
XP12Bb  B12  B12B  INV
XP13Bb  B13  B13B  INV
XP14Bb  B14  B14B  INV
XP15Bb  B15  B15B  INV
XP16Bb  B16  B16B  INV
XP17Bb  B17  B17B  INV
XP18Bb  B18  B18B  INV
XP19Bb  B19  B19B  INV
XP20Bb  B20  B20B  INV
XP21Bb  B21  B21B  INV
XP22Bb  B22  B22B  INV
XP23Bb  B23  B23B  INV
XP24Bb  B24  B24B  INV
XP25Bb  B25  B25B  INV
XP26Bb  B26  B26B  INV
XP27Bb  B27  B27B  INV
XP28Bb  B28  B28B  INV
XP29Bb  B29  B29B  INV
XP30Bb  B30  B30B  INV
XP31Bb  B31  B31B  INV
      ********************Inverse P**********
XP0Pb  P0  P0B  INV   M='HINV' 
XP1Pb  P1  P1B  INV   M='HINV'
XP2Pb  P2  P2B  INV   M='HINV'
XP3Pb  P3  P3B  INV   M='HINV'
XP4Pb  P4  P4B  INV   M='HINV'
XP5Pb  P5  P5B  INV   M='HINV'
XP6Pb  P6  P6B  INV   M='HINV'
XP7Pb  P7  P7B  INV   M='HINV'
XP8Pb  P8  P8B  INV   M='HINV'
XP9Pb  P9  P9B  INV   M='HINV'
XP10Pb  P10  P10B  INV   M='HINV'  
XP11Pb  P11  P11B  INV   M='HINV'
XP12Pb  P12  P12B  INV   M='HINV'
XP13Pb  P13  P13B  INV   M='HINV'
XP14Pb  P14  P14B  INV   M='HINV'
XP15Pb  P15  P15B  INV   M='HINV'
XP16Pb  P16  P16B  INV   M='HINV'
XP17Pb  P17  P17B  INV   M='HINV'
XP18Pb  P18  P18B  INV   M='HINV'
XP19Pb  P19  P19B  INV   M='HINV'
XP20Pb  P20  P20B  INV   M='HINV'
XP21Pb  P21  P21B  INV   M='HINV'
XP22Pb  P22  P22B  INV   M='HINV'
XP23Pb  P23  P23B  INV   M='HINV'
XP24Pb  P24  P24B  INV   M='HINV'
XP25Pb  P25  P25B  INV   M='HINV'
XP26Pb  P26  P26B  INV   M='HINV'
XP27Pb  P27  P27B  INV   M='HINV'
XP28Pb  P28  P28B  INV   M='HINV'
XP29Pb  P29  P29B  INV   M='HINV'
XP30Pb  P30  P30B  INV   M='HINV'
XP31Pb  P31  P31B  INV   M='HINV'

***********Propagate 1st Level**************
XP0  A0  B0  A0B   B0B   CLK   P0   PROP   M='H1'
XP1  A1  B1  A1B   B1B   CLK   P1   PROP   M='H1'
XP2  A2  B2  A2B   B2B   CLK   P2   PROP   M='H1'
XP3  A3  B3  A3B   B3B   CLK   P3   PROP   M='H1'
XP4  A4  B4  A4B   B4B   CLK   P4   PROP   M='H1'
XP5  A5  B5  A5B   B5B   CLK   P5   PROP   M='H1'
XP6  A6  B6  A6B   B6B   CLK   P6   PROP   M='H1'
XP7  A7  B7  A7B   B7B   CLK   P7   PROP   M='H1'
XP8  A8  B8  A8B   B8B   CLK   P8   PROP   M='H1'
XP9  A9  B9  A9B   B9B   CLK   P9   PROP   M='H1'
XP10   A10   B10   A10B   B10B CLK P10   PROP   M='H1'
XP11   A11   B11   A11B   B11B CLK P11   PROP   M='H1'
XP12   A12   B12   A12B   B12B CLK P12   PROP   M='H1'
XP13   A13   B13   A13B   B13B CLK P13   PROP   M='H1'
XP14   A14   B14   A14B   B14B CLK P14   PROP   M='H1'
XP15   A15   B15   A15B   B15B CLK P15   PROP   M='H1'
XP16   A16   B16   A16B   B16B CLK P16   PROP   M='H1'
XP17   A17   B17   A17B   B17B CLK P17   PROP   M='H1'
XP18   A18   B18   A18B   B18B CLK P18   PROP   M='H1'
XP19   A19   B19   A19B   B19B CLK P19   PROP   M='H1'
XP20   A20   B20   A20B   B20B CLK P20   PROP   M='H1'
XP21   A21   B21   A21B   B21B CLK P21   PROP   M='H1'
XP22   A22   B22   A22B   B22B CLK P22   PROP   M='H1'
XP23   A23   B23   A23B   B23B CLK P23   PROP   M='H1'
XP24   A24   B24   A24B   B24B CLK P24   PROP   M='H1'
XP25   A25   B25   A25B   B25B CLK P25   PROP   M='H1'
XP26   A26   B26   A26B   B26B CLK P26   PROP   M='H1'
XP27   A27   B27   A27B   B27B CLK P27   PROP   M='H1'
XP28   A28   B28   A28B   B28B CLK P28   PROP   M='H1'
XP29   A29   B29   A29B   B29B CLK P29   PROP   M='H1'
XP30   A30   B30   A30B   B30B CLK P30   PROP   M='H1'
XP31   A31   B31   A31B   B31B CLK P31   PROP   M='H1'
  
***********Generate 1st Level**************
XG0  A0  B0  CLK  G0  GENERATE  M='H2'
XG1  A1  B1  CLK  G1  GENERATE  M='H2'
XG2  A2  B2  CLK  G2  GENERATE  M='H2'
XG3  A3  B3  CLK  G3  GENERATE  M='H2'
XG4  A4  B4  CLK  G4  GENERATE  M='H2'
XG5  A5  B5  CLK  G5  GENERATE  M='H2'
XG6  A6  B6  CLK  G6  GENERATE  M='H2'
XG7  A7  B7  CLK  G7  GENERATE  M='H2'
XG8  A8  B8  CLK  G8  GENERATE  M='H2'
XG9  A9  B9  CLK  G9  GENERATE  M='H2'
XG10  A10  B10  CLK  G10  GENERATE  M='H2'
XG11  A11  B11  CLK  G11  GENERATE  M='H2'
XG12  A12  B12  CLK  G12  GENERATE  M='H2'
XG13  A13  B13  CLK  G13  GENERATE  M='H2'
XG14  A14  B14  CLK  G14  GENERATE  M='H2'
XG15  A15  B15  CLK  G15  GENERATE  M='H2'
XG16  A16  B16  CLK  G16  GENERATE  M='H2'
XG17  A17  B17  CLK  G17  GENERATE  M='H2'
XG18  A18  B18  CLK  G18  GENERATE  M='H2'
XG19  A19  B19  CLK  G19  GENERATE  M='H2'
XG20  A20  B20  CLK  G20  GENERATE  M='H2'
XG21  A21  B21  CLK  G21  GENERATE  M='H2'
XG22  A22  B22  CLK  G22  GENERATE  M='H2'
XG23  A23  B23  CLK  G23  GENERATE  M='H2'
XG24  A24  B24  CLK  G24  GENERATE  M='H2'
XG25  A25  B25  CLK  G25  GENERATE  M='H2'
XG26  A26  B26  CLK  G26  GENERATE  M='H2'
XG27  A27  B27  CLK  G27  GENERATE  M='H2'
XG28  A28  B28  CLK  G28  GENERATE  M='H2'
XG29  A29  B29  CLK  G29  GENERATE  M='H2'
XG30  A30  B30  CLK  G30  GENERATE  M='H2'
XG31  A31  B31  CLK  G31  GENERATE  M='H2'
***********DOT 1st Level(Level: 32-1=31)**************
XDOT1_0   G0  P0  G1  P1  G1_0   P1_0	CLK  DOT   M='H3'
XDOT1_1   G1  P1  G2  P2  G2_1   P2_1	CLK  DOT   M='H3'
XDOT1_2   G2  P2  G3  P3  G3_2   P3_2	CLK  DOT   M='H3'
XDOT1_3   G3  P3  G4  P4  G4_3   P4_3	CLK  DOT   M='H3'
XDOT1_4   G4  P4  G5  P5  G5_4   P5_4	CLK  DOT   M='H3'
XDOT1_5   G5  P5  G6  P6  G6_5   P6_5	CLK  DOT   M='H3'
XDOT1_6   G6  P6  G7  P7  G7_6   P7_6	CLK  DOT   M='H3'
XDOT1_7   G7  P7  G8  P8  G8_7   P8_7	CLK  DOT   M='H3'
XDOT1_8   G8  P8  G9  P9  G9_8   P9_8	CLK  DOT   M='H3'
XDOT1_9   G9  P9  G10 P10  G10_9   P10_9 CLK  DOT   M='H3'
XDOT1_10  G10  P10  G11  P11  G11_10   P11_10 CLK  DOT   M='H3'
XDOT1_11  G11  P11  G12  P12  G12_11   P12_11 CLK  DOT   M='H3'
XDOT1_12  G12  P12  G13  P13  G13_12   P13_12 CLK  DOT   M='H3'
XDOT1_13  G13  P13  G14  P14  G14_13   P14_13 CLK  DOT   M='H3'
XDOT1_14  G14  P14  G15  P15  G15_14   P15_14 CLK  DOT   M='H3'
XDOT1_15  G15  P15  G16  P16  G16_15   P16_15 CLK  DOT   M='H3'
XDOT1_16  G16  P16  G17  P17  G17_16   P17_16 CLK  DOT   M='H3'
XDOT1_17  G17  P17  G18  P18  G18_17   P18_17 CLK  DOT   M='H3'
XDOT1_18  G18  P18  G19  P19  G19_18   P19_18 CLK  DOT   M='H3'
XDOT1_19  G19  P19  G20  P20  G20_19   P20_19 CLK  DOT   M='H3'
XDOT1_20  G20  P20  G21  P21  G21_20   P21_20 CLK  DOT   M='H3'
XDOT1_21  G21  P21  G22  P22  G22_21   P22_21 CLK  DOT   M='H3'
XDOT1_22  G22  P22  G23  P23  G23_22   P23_22 CLK  DOT   M='H3'
XDOT1_23  G23  P23  G24  P24  G24_23   P24_23 CLK  DOT   M='H3'
XDOT1_24  G24  P24  G25  P25  G25_24   P25_24 CLK  DOT   M='H3'
XDOT1_25  G25  P25  G26  P26  G26_25   P26_25 CLK  DOT   M='H3'
XDOT1_26  G26  P26  G27  P27  G27_26   P27_26 CLK  DOT   M='H3'
XDOT1_27  G27  P27  G28  P28  G28_27   P28_27 CLK  DOT   M='H3'
XDOT1_28  G28  P28  G29  P29  G29_28   P29_28 CLK  DOT   M='H3'
XDOT1_29  G29  P29  G30  P30  G30_29   P30_29 CLK  DOT   M='H3'
XDOT1_30  G30  P30  G31  P31  G31_30   P31_30 CLK  DOT   M='H3'

***********DOT 2nd Level(Level: 32-2=30)**************
XDOT2_0  G0     P0      G2_1    P2_1    G2_0    P2_0   CLK  DOT   M='H4'
XDOT2_1  G1_0   P1_0    G3_2    P3_2    G3_0    P3_0   CLK  DOT   M='H4'
XDOT2_2  G2_1   P2_1    G4_3    P4_3    G4_1    P4_1   CLK  DOT   M='H4'
XDOT2_3  G3_2   P3_2    G5_4    P5_4    G5_2    P5_2   CLK  DOT   M='H4'
XDOT2_4  G4_3   P4_3    G6_5    P6_5    G6_3    P6_3   CLK  DOT   M='H4'
XDOT2_5  G5_4   P5_4    G7_6    P7_6    G7_4    P7_4   CLK  DOT   M='H4'
XDOT2_6  G6_5   P6_5    G8_7    P8_7    G8_5    P8_5   CLK  DOT   M='H4'
XDOT2_7  G7_6   P7_6    G9_8    P9_8    G9_6    P9_6   CLK  DOT   M='H4'
XDOT2_8  G8_7   P8_7    G10_9   P10_9   G10_7   P10_7  CLK  DOT   M='H4'
XDOT2_9  G9_8   P9_8    G11_10  P11_10  G11_8   P11_8  CLK  DOT   M='H4'
XDOT2_10  G10_9  P10_9  G12_11  P12_11  G12_9   P12_9  CLK  DOT	M='H4'
XDOT2_11  G11_10   P11_10	G13_12	P13_12	G13_10	P13_10	CLK  DOT	M='H4'
XDOT2_12  G12_11   P12_11	G14_13	P14_13	G14_11	P14_11	CLK  DOT	M='H4'
XDOT2_13  G13_12   P13_12	G15_14	P15_14	G15_12	P15_12	CLK  DOT	M='H4'
XDOT2_14  G14_13   P14_13	G16_15	P16_15	G16_13	P16_13	CLK  DOT	M='H4'
XDOT2_15  G15_14   P15_14	G17_16	P17_16	G17_14	P17_14	CLK  DOT	M='H4'
XDOT2_16  G16_15   P16_15	G18_17	P18_17	G18_15	P18_15	CLK  DOT	M='H4'
XDOT2_17  G17_16   P17_16	G19_18	P19_18	G19_16	P19_16	CLK  DOT	M='H4'
XDOT2_18  G18_17   P18_17	G20_19	P20_19	G20_17	P20_17	CLK  DOT	M='H4'
XDOT2_19  G19_18   P19_18	G21_20	P21_20	G21_18	P21_18	CLK  DOT	M='H4'
XDOT2_20  G20_19   P20_19	G22_21	P22_21	G22_19	P22_19	CLK  DOT	M='H4'
XDOT2_21  G21_20   P21_20	G23_22	P23_22	G23_20	P23_20	CLK  DOT	M='H4'
XDOT2_22  G22_21   P22_21	G24_23	P24_23	G24_21	P24_21	CLK  DOT	M='H4'
XDOT2_23  G23_22   P23_22	G25_24	P25_24	G25_22	P25_22	CLK  DOT	M='H4'
XDOT2_24  G24_23   P24_23	G26_25	P26_25	G26_23	P26_23	CLK  DOT	M='H4'
XDOT2_25  G25_24   P25_24	G27_26	P27_26	G27_24	P27_24	CLK  DOT	M='H4'
XDOT2_26  G26_25   P26_25	G28_27	P28_27	G28_25	P28_25	CLK  DOT	M='H4'
XDOT2_27  G27_26   P27_26	G29_28	P29_28	G29_26	P29_26	CLK  DOT	M='H4'
XDOT2_28  G28_27   P28_27	G30_29	P30_29	G30_27	P30_27	CLK  DOT	M='H4'
XDOT2_29  G29_28   P29_28	G31_30	P31_30	G31_28	P31_28	CLK  DOT	M='H4'

***********DOT 3rd Level(Level: 32-4=28)**************
XDOT3_0     G0	    P0	G4_1	P4_1	G4_0	P4_0	CLK DOT	M='H5'
XDOT3_1     G1_0	P1_0	G5_2	P5_2	G5_0	P5_0	CLK  DOT	M='H5'
XDOT3_2     G2_0	P2_0	G6_3	P6_3	G6_0	P6_0	CLK  DOT	M='H5'
XDOT3_3     G3_0	P3_0	G7_4	P7_4	G7_0	P7_0	CLK  DOT	M='H5'
XDOT3_4     G4_1	P4_1	G8_5	P8_5	G8_1	P8_1	CLK  DOT	M='H5'
XDOT3_5     G5_2	P5_2	G9_6	P9_6	G9_2	P9_2	CLK  DOT	M='H5'
XDOT3_6     G6_3	P6_3	G10_7	P10_7	G10_3	P10_3	CLK  DOT	M='H5'
XDOT3_7     G7_4	P7_4	G11_8	P11_8	G11_4	P11_4	CLK  DOT	M='H5'
XDOT3_8     G8_5	P8_5	G12_9	P12_9	G12_5	P12_5	CLK  DOT	M='H5'
XDOT3_9		G9_6	P9_6	G13_10	P13_10	G13_6	P13_6	CLK  DOT	M='H5'
XDOT3_10	G10_7	P10_7	G14_11	P14_11	G14_7	P14_7	CLK  DOT	M='H5'
XDOT3_11	G11_8	P11_8	G15_12	P15_12	G15_8	P15_8	CLK  DOT	M='H5'
XDOT3_12	G12_9	P12_9	G16_13	P16_13	G16_9	P16_9	CLK  DOT	M='H5'
XDOT3_13	G13_10	P13_10	G17_14	P17_14	G17_10	P17_10	CLK  DOT	M='H5'
XDOT3_14	G14_11	P14_11	G18_15	P18_15	G18_11	P18_11	CLK  DOT	M='H5'
XDOT3_15	G15_12	P15_12	G19_16	P19_16	G19_12	P19_12	CLK  DOT	M='H5'
XDOT3_16	G16_13	P16_13	G20_17	P20_17	G20_13	P20_13	CLK  DOT	M='H5'
XDOT3_17	G17_14	P17_14	G21_18	P21_18	G21_14	P21_14	CLK  DOT	M='H5'
XDOT3_18	G18_15	P18_15	G22_19	P22_19	G22_15	P22_15	CLK  DOT	M='H5'
XDOT3_19	G19_16	P19_16	G23_20	P23_20	G23_16	P23_16	CLK  DOT	M='H5'
XDOT3_20	G20_17	P20_17	G24_21	P24_21	G24_17	P24_17	CLK  DOT	M='H5'
XDOT3_21	G21_18	P21_18	G25_22	P25_22	G25_18	P25_18	CLK  DOT	M='H5'
XDOT3_22	G22_19	P22_19	G26_23	P26_23	G26_19	P26_19	CLK  DOT	M='H5'
XDOT3_23	G23_20	P23_20	G27_24	P27_24	G27_20	P27_20	CLK  DOT	M='H5'
XDOT3_24	G24_21	P24_21	G28_25	P28_25	G28_21	P28_21	CLK  DOT	M='H5'
XDOT3_25	G25_22	P25_22	G29_26	P29_26	G29_22	P29_22	CLK  DOT	M='H5'
XDOT3_26	G26_23	P26_23	G30_27	P30_27	G30_23	P30_23	CLK  DOT	M='H5'
XDOT3_27	G27_24	P27_24	G31_28	P31_28	G31_24	P31_24	CLK  DOT	M='H5'

***********DOT 4th Level(Level: 32-8=24)**************
XDOT4_0  G0	P0	G8_1	P8_1	G8_0	P8_0	CLK  DOT	M='H6'
XDOT4_1  G1_0	P1_0	G9_2	P9_2	G9_0	P9_0	CLK  DOT	M='H6'
XDOT4_2  G2_0	P2_0	G10_3	P10_3	G10_0	P10_0	CLK  DOT	M='H6'
XDOT4_3  G3_0	P3_0	G11_4	P11_4	G11_0	P11_0	CLK  DOT	M='H6'
XDOT4_4  G4_0	P4_0	G12_5	P12_5	G12_0	P12_0	CLK  DOT	M='H6'
XDOT4_5  G5_0	P5_0	G13_6	P13_6	G13_0	P13_0	CLK  DOT	M='H6'
XDOT4_6  G6_0	P6_0	G14_7	P14_7	G14_0	P14_0	CLK  DOT	M='H6'
XDOT4_7  G7_0	P7_0	G15_8	P15_8	G15_0	P15_0	CLK  DOT	M='H6'
XDOT4_8  G8_1	P8_1	G16_9	P16_9	G16_1	P16_1	CLK  DOT	M='H6'
XDOT4_9  G9_2	P9_2	G17_10	P17_10	G17_2	P17_2	CLK  DOT	M='H6'
XDOT4_10 G10_3	P10_3	G18_11	P18_11	G18_3	P18_3	CLK  DOT	M='H6'
XDOT4_11 G11_4	P11_4	G19_12	P19_12	G19_4	P19_4	CLK  DOT	M='H6'
XDOT4_12 G12_5	P12_5	G20_13	P20_13	G20_5	P20_5	CLK  DOT	M='H6'
XDOT4_13 G13_6	P13_6	G21_14	P21_14	G21_6	P21_6	CLK  DOT	M='H6'
XDOT4_14 G14_7	P14_7	G22_15	P22_15	G22_7	P22_7	CLK  DOT	M='H6'
XDOT4_15 G15_8	P15_8	G23_16	P23_16	G23_8	P23_8	CLK  DOT	M='H6'
XDOT4_16 G16_9	P16_9	G24_17	P24_17	G24_9	P24_9	CLK  DOT	M='H6'
XDOT4_17 G17_10	P17_10	G25_18	P25_18	G25_10	P25_10	CLK  DOT	M='H6'
XDOT4_18 G18_11	P18_11	G26_19	P26_19	G26_11	P26_11	CLK  DOT	M='H6'
XDOT4_19 G19_12	P19_12	G27_20	P27_20	G27_12	P27_12	CLK  DOT	M='H6'
XDOT4_20 G20_13	P20_13	G28_21	P28_21	G28_13	P28_13	CLK  DOT	M='H6'
XDOT4_21 G21_14	P21_14	G29_22	P29_22	G29_14	P29_14	CLK  DOT	M='H6'
XDOT4_22 G22_15	P22_15	G30_23	P30_23	G30_15	P30_15	CLK  DOT	M='H6'
XDOT4_23 G23_16	P23_16	G31_24	P31_24	G31_16	P31_16	CLK  DOT	M='H6'

***********DOT 5th Level(Level: 32-16=16)**************
XODT5_0    G0       P0      G16_1   P16_1	G16_0	P16_0	CLK  DOT	M='H7'
XDOT5_1    G1_0     P1_0    G17_2   P17_2	G17_0	P17_0	CLK  DOT	M='H7'
XDOT5_2    G2_0     P2_0    G18_3   P18_3	G18_0	P18_0	CLK  DOT	M='H7'
XDOT5_3    G3_0     P3_0    G19_4   P19_4	G19_0	P19_0	CLK  DOT	M='H7'
XDOT5_4    G4_0     P4_0    G20_5   P20_5	G20_0	P20_0	CLK  DOT	M='H7'
XDOT5_5    G5_0     P5_0    G21_6   P21_6	G21_0	P21_0	CLK  DOT	M='H7'
XDOT5_6    G6_0     P6_0    G22_7   P22_7	G22_0	P22_0	CLK  DOT	M='H7'
XDOT5_7    G7_0     P7_0    G23_8   P23_8	G23_0	P23_0	CLK  DOT	M='H7'
XDOT5_8    G8_0     P8_0    G24_9   P24_9	G24_0	P24_0	CLK  DOT	M='H7'
XDOT5_9    G9_0     P9_0    G25_10  P25_10	G25_0	P25_0	CLK  DOT	M='H7'
XDOT5_10   G10_0    P10_0   G26_11  P26_11	G26_0	P26_0	CLK  DOT	M='H7'
XDOT5_11   G11_0    P11_0   G27_12  P27_12	G27_0	P27_0	CLK  DOT	M='H7'
XDOT5_12   G12_0    P12_0   G28_13  P28_13	G28_0	P28_0	CLK  DOT	M='H7'
XDOT5_13   G13_0    P13_0   G29_14  P29_14	G29_0	P29_0	CLK  DOT	M='H7'
XDOT5_14   G14_0    P14_0   G30_15  P30_15	G30_0	P30_0	CLK  DOT	M='H7'
XDOT5_15   G15_0    P15_0   G31_16  P31_16	G31_0	P31_0	CLK  DOT	M='H7'

***********SUM**************
XSUM0	P0	P0B  GND	CLK  CLK_D  S0	SUM   M='H8'
XSUM1	P1	P1B  G0	    CLK  CLK_D  S1	SUM   M='H8'
XSUM2	P2	P2B  G1_0	CLK  CLK_D  S2	SUM   M='H8'
XSUM3	P3	P3B  G2_0	CLK  CLK_D  S3	SUM   M='H8'
XSUM4	P4	P4B  G3_0	CLK  CLK_D  S4	SUM   M='H8'
XSUM5	P5	P5B  G4_0	CLK  CLK_D  S5	SUM   M='H8'
XSUM6	P6	P6B  G5_0	CLK  CLK_D  S6	SUM   M='H8'
XSUM7	P7	P7B  G6_0	CLK  CLK_D  S7	SUM   M='H8'
XSUM8	P8	P8B  G7_0	CLK  CLK_D  S8	SUM   M='H8'
XSUM9	P9	P9B  G8_0	CLK  CLK_D  S9	SUM   M='H8'
XSUM10	P10	P10B G9_0	CLK  CLK_D  S10	SUM   M='H8'
XSUM11	P11	P11B G10_0	CLK  CLK_D  S11	SUM   M='H8'
XSUM12	P12	P12B G11_0	CLK  CLK_D  S12	SUM   M='H8'
XSUM13	P13	P13B G12_0	CLK  CLK_D  S13	SUM   M='H8'
XSUM14	P14	P14B G13_0	CLK  CLK_D  S14	SUM   M='H8'
XSUM15	P15	P15B G14_0	CLK  CLK_D  S15	SUM   M='H8'
XSUM16	P16	P16B G15_0	CLK  CLK_D  S16	SUM   M='H8'
XSUM17	P17	P17B G16_0	CLK  CLK_D  S17	SUM   M='H8'
XSUM18	P18	P18B G17_0	CLK  CLK_D  S18	SUM   M='H8'
XSUM19	P19	P19B G18_0	CLK  CLK_D  S19	SUM   M='H8'
XSUM20	P20	P20B G19_0	CLK  CLK_D  S20	SUM   M='H8'
XSUM21	P21	P21B G20_0	CLK  CLK_D  S21	SUM   M='H8'
XSUM22	P22	P22B G21_0	CLK  CLK_D  S22	SUM   M='H8'
XSUM23	P23	P23B G22_0	CLK  CLK_D  S23	SUM   M='H8'
XSUM24	P24	P24B G23_0	CLK  CLK_D  S24	SUM   M='H8'
XSUM25	P25	P25B G24_0	CLK  CLK_D  S25	SUM   M='H8'
XSUM26	P26	P26B G25_0	CLK  CLK_D  S26	SUM   M='H8'
XSUM27	P27	P27B G26_0	CLK  CLK_D  S27	SUM   M='H8'
XSUM28	P28	P28B G27_0	CLK  CLK_D  S28	SUM   M='H8'
XSUM29	P29	P29B G28_0	CLK  CLK_D  S29	SUM   M='H8'
XSUM30	P30	P30B G29_0	CLK  CLK_D  S30	SUM   M='H8'
XSUM31	P31	P31B G30_0	CLK  CLK_D  S31	SUM   M='H8'


**********************Source*****************
VDD VDD GND '0.85'
VCLK CLK GND PULSE 0 'SUPPLY' 50ps 15ps 15ps 470ps 1ns
VCLK_D CLK_D GND PULSE 0 'SUPPLY' 59ps 15ps 15ps 470ps 1ns

.vec lp_stimulus.vect
.tran 1ps 8ns 
.op all 
.measure TRAN leakage_power AVG P(VDD) FROM=0ns TO=8ns
.end