.TITLE ADDER
.lib "..\models" ptm16lstp
.options acct list post
.global vdd gnd vss vdda
.TEMP 85

.param D=1
.param H=1
.param vds_sup=0.1
.param supply=0.85

.param finp=1
.param finn=1
.param length=20n
.param fint=12n
.param finh=26n

.param L1=1
.param L2=2
.param L3=3
.param L4=4
.param L5=5
.param L6=6
.param L7=7
.param L8=8
*
.SUBCKT INV A Y nfinn=finn nfinp=finp
xnmos Y A GND GND lnfet l=length nfin=nfinn
xpmos Y A VDD VDD lpfet l=length nfin=nfinp
.ENDS
*
.SUBCKT XOR2 A B P nfinn=finn nfinp=finp
* generate signal P
xpmos1 N1 B VDD VDD lpfet l=length nfin=nfinp 
xpmos2 X1 A N1 VDD lpfet l=length nfin=nfinp 
xpmos3 N2 B VDD VDD lpfet l=length nfin=nfinp 
xpmos4 N2 A VDD VDD lpfet l=length nfin=nfinp 
xpmos5 P X1 N2 VDD lpfet l=length nfin=nfinp 

xnmos1 X1 B GND GND lnfet l=length nfin=nfinn
xnmos2 X1 A GND GND lnfet l=length nfin=nfinn
xnmos3 P A N3 GND lnfet l=length nfin=nfinn
xnmos4 N3 B GND GND lnfet l=length nfin=nfinn
xnmos5 P X1 GND GND lnfet l=length nfin=nfinn
.ENDS

.SUBCKT AND2 A B G nfinn=finn nfinp=finp
* generate signal G
xpmos6 X2 A VDD VDD lpfet l=length nfin=nfinp 
xpmos7 X2 B VDD VDD lpfet l=length nfin=nfinp 
xpmos8 G X2 VDD VDD lpfet l=length nfin=nfinp 

xnmos6 X2 B N4 GND lnfet l=length nfin=nfinn
xnmos7 N4 A GND GND lnfet l=length nfin=nfinn
xnmos8 G X2 GND GND lnfet l=length nfin=nfinn

.ENDS
*
.SUBCKT OR2 A B Y nfinn=finn nfinp=finp
xpmos9 N5 A VDD VDD lpfet l=length nfin=nfinp 
xpmos10 X3 B N5 VDD lpfet l=length nfin=nfinp 
xpmos11 Y X3 VDD VDD lpfet l=length nfin=nfinp 

xnmos9 X3 A GND GND lnfet l=length nfin=nfinn
xnmos10 X3 B GND GND lnfet l=length nfin=nfinn
xnmos11 Y X3 GND GND lnfet l=length nfin=nfinn

.ENDS

.SUBCKT DOT G1 P1 G2 P2 GOUT POUT D=H
XAND1 P1 G2 P1G2 AND2 M='H'
XOR1 G1 P1G2 GOUT OR2 M='H'
XAND2 P1 P2 POUT AND2 M='H'
.ENDS

*P generation
XP0	A0	B0	P0	XOR2	M='L1'
XP1	A1	B1	P1	XOR2	M='L1'
XP2	A2	B2	P2	XOR2	M='L1'
XP3	A3	B3	P3	XOR2	M='L1'
XP4	A4	B4	P4	XOR2	M='L1'
XP5	A5	B5	P5	XOR2	M='L1'
XP6	A6	B6	P6	XOR2	M='L1'
XP7	A7	B7	P7	XOR2	M='L1'
XP8	A8	B8	P8	XOR2	M='L1'
XP9	A9	B9	P9	XOR2	M='L1'
XP10	A10	B10	P10	XOR2	M='L1'
XP11	A11	B11	P11	XOR2	M='L1'
XP12	A12	B12	P12	XOR2	M='L1'
XP13	A13	B13	P13	XOR2	M='L1'
XP14	A14	B14	P14	XOR2	M='L1'
XP15	A15	B15	P15	XOR2	M='L1'
XP16	A16	B16	P16	XOR2	M='L1'
XP17	A17	B17	P17	XOR2	M='L1'
XP18	A18	B18	P18	XOR2	M='L1'
XP19	A19	B19	P19	XOR2	M='L1'
XP20	A20	B20	P20	XOR2	M='L1'
XP21	A21	B21	P21	XOR2	M='L1'
XP22	A22	B22	P22	XOR2	M='L1'
XP23	A23	B23	P23	XOR2	M='L1'
XP24	A24	B24	P24	XOR2	M='L1'
XP25	A25	B25	P25	XOR2	M='L1'
XP26	A26	B26	P26	XOR2	M='L1'
XP27	A27	B27	P27	XOR2	M='L1'
XP28	A28	B28	P28	XOR2	M='L1'
XP29	A29	B29	P29	XOR2	M='L1'
XP30	A30	B30	P30	XOR2	M='L1'
XP31	A31	B31	P31	XOR2	M='L1'

*P generation
XG0	A0	B0	G0	AND2	M='L2'
XG1	A1	B1	G1	AND2	M='L2'
XG2	A2	B2	G2	AND2	M='L2'
XG3	A3	B3	G3	AND2	M='L2'
XG4	A4	B4	G4	AND2	M='L2'
XG5	A5	B5	G5	AND2	M='L2'
XG6	A6	B6	G6	AND2	M='L2'
XG7	A7	B7	G7	AND2	M='L2'
XG8	A8	B8	G8	AND2	M='L2'
XG9	A9	B9	G9	AND2	M='L2'
XG10	A10	B10	G10	AND2	M='L2'
XG11	A11	B11	G11	AND2	M='L2'
XG12	A12	B12	G12	AND2	M='L2'
XG13	A13	B13	G13	AND2	M='L2'
XG14	A14	B14	G14	AND2	M='L2'
XG15	A15	B15	G15	AND2	M='L2'
XG16	A16	B16	G16	AND2	M='L2'
XG17	A17	B17	G17	AND2	M='L2'
XG18	A18	B18	G18	AND2	M='L2'
XG19	A19	B19	G19	AND2	M='L2'
XG20	A20	B20	G20	AND2	M='L2'
XG21	A21	B21	G21	AND2	M='L2'
XG22	A22	B22	G22	AND2	M='L2'
XG23	A23	B23	G23	AND2	M='L2'
XG24	A24	B24	G24	AND2	M='L2'
XG25	A25	B25	G25	AND2	M='L2'
XG26	A26	B26	G26	AND2	M='L2'
XG27	A27	B27	G27	AND2	M='L2'
XG28	A28	B28	G28	AND2	M='L2'
XG29	A29	B29	G29	AND2	M='L2'
XG30	A30	B30	G30	AND2	M='L2'
XG31	A31	B31	G31	AND2	M='L2'

XDOT0	G0	P0	G1	P1	G1_0	P1_0	DOT	M='L3'
XDOT1	G1	P1	G2	P2	G2_1	P2_1	DOT	M='L3'
XDOT2	G2	P2	G3	P3	G3_2	P3_2	DOT	M='L3'
XDOT3	G3	P3	G4	P4	G4_3	P4_3	DOT	M='L3'
XDOT4	G4	P4	G5	P5	G5_4	P5_4	DOT	M='L3'
XDOT5	G5	P5	G6	P6	G6_5	P6_5	DOT	M='L3'
XDOT6	G6	P6	G7	P7	G7_6	P7_6	DOT	M='L3'
XDOT7	G7	P7	G8	P8	G8_7	P8_7	DOT	M='L3'
XDOT8	G8	P8	G9	P9	G9_8	P9_8	DOT	M='L3'
XDOT9	G9	P9	G10	P10	G10_9	P10_9	DOT	M='L3'
XDOT10	G10	P10	G11	P11	G11_10	P11_10	DOT	M='L3'
XDOT11	G11	P11	G12	P12	G12_11	P12_11	DOT	M='L3'
XDOT12	G12	P12	G13	P13	G13_12	P13_12	DOT	M='L3'
XDOT13	G13	P13	G14	P14	G14_13	P14_13	DOT	M='L3'
XDOT14	G14	P14	G15	P15	G15_14	P15_14	DOT	M='L3'
XDOT15	G15	P15	G16	P16	G16_15	P16_15	DOT	M='L3'
XDOT16	G16	P16	G17	P17	G17_16	P17_16	DOT	M='L3'
XDOT17	G17	P17	G18	P18	G18_17	P18_17	DOT	M='L3'
XDOT18	G18	P18	G19	P19	G19_18	P19_18	DOT	M='L3'
XDOT19	G19	P19	G20	P20	G20_19	P20_19	DOT	M='L3'
XDOT20	G20	P20	G21	P21	G21_20	P21_20	DOT	M='L3'
XDOT21	G21	P21	G22	P22	G22_21	P22_21	DOT	M='L3'
XDOT22	G22	P22	G23	P23	G23_22	P23_22	DOT	M='L3'
XDOT23	G23	P23	G24	P24	G24_23	P24_23	DOT	M='L3'
XDOT24	G24	P24	G25	P25	G25_24	P25_24	DOT	M='L3'
XDOT25	G25	P25	G26	P26	G26_25	P26_25	DOT	M='L3'
XDOT26	G26	P26	G27	P27	G27_26	P27_26	DOT	M='L3'
XDOT27	G27	P27	G28	P28	G28_27	P28_27	DOT	M='L3'
XDOT28	G28	P28	G29	P29	G29_28	P29_28	DOT	M='L3'
XDOT29	G29	P29	G30	P30	G30_29	P30_29	DOT	M='L3'
XDOT30	G30	P30	G31	P31	G31_30	P31_30	DOT	M='L3'

*level 2 signal
XDOT31	G0	P0	G2_1	P2_1	G2_0	P2_0	DOT	M='L4'
XDOT32	G1_0	P1_0	G3_2	P3_2	G3_0	P3_0	DOT	M='L4'
XDOT33	G2_1	P2_1	G4_3	P4_3	G4_1	P4_1	DOT	M='L4'
XDOT34	G3_2	P3_2	G5_4	P5_4	G5_2	P5_2	DOT	M='L4'
XDOT35	G4_3	P4_3	G6_5	P6_5	G6_3	P6_3	DOT	M='L4'
XDOT36	G5_4	P5_4	G7_6	P7_6	G7_4	P7_4	DOT	M='L4'
XDOT37	G6_5	P6_5	G8_7	P8_7	G8_5	P8_5	DOT	M='L4'
XDOT38	G7_6	P7_6	G9_8	P9_8	G9_6	P9_6	DOT	M='L4'
XDOT39	G8_7	P8_7	G10_9	P10_9	G10_7	P10_7	DOT	M='L4'
XDOT40	G9_8	P9_8	G11_10	P11_10	G11_8	P11_8	DOT	M='L4'
XDOT41	G10_9	P10_9	G12_11	P12_11	G12_9	P12_9	DOT	M='L4'
XDOT42	G11_10	P11_10	G13_12	P13_12	G13_10	P13_10	DOT	M='L4'
XDOT43	G12_11	P12_11	G14_13	P14_13	G14_11	P14_11	DOT	M='L4'
XDOT44	G13_12	P13_12	G15_14	P15_14	G15_12	P15_12	DOT	M='L4'
XDOT45	G14_13	P14_13	G16_15	P16_15	G16_13	P16_13	DOT	M='L4'
XDOT46	G15_14	P15_14	G17_16	P17_16	G17_14	P17_14	DOT	M='L4'
XDOT47	G16_15	P16_15	G18_17	P18_17	G18_15	P18_15	DOT	M='L4'
XDOT48	G17_16	P17_16	G19_18	P19_18	G19_16	P19_16	DOT	M='L4'
XDOT49	G18_17	P18_17	G20_19	P20_19	G20_17	P20_17	DOT	M='L4'
XDOT50	G19_18	P19_18	G21_20	P21_20	G21_18	P21_18	DOT	M='L4'
XDOT51	G20_19	P20_19	G22_21	P22_21	G22_19	P22_19	DOT	M='L4'
XDOT52	G21_20	P21_20	G23_22	P23_22	G23_20	P23_20	DOT	M='L4'
XDOT53	G22_21	P22_21	G24_23	P24_23	G24_21	P24_21	DOT	M='L4'
XDOT54	G23_22	P23_22	G25_24	P25_24	G25_22	P25_22	DOT	M='L4'
XDOT55	G24_23	P24_23	G26_25	P26_25	G26_23	P26_23	DOT	M='L4'
XDOT56	G25_24	P25_24	G27_26	P27_26	G27_24	P27_24	DOT	M='L4'
XDOT57	G26_25	P26_25	G28_27	P28_27	G28_25	P28_25	DOT	M='L4'
XDOT58	G27_26	P27_26	G29_28	P29_28	G29_26	P29_26	DOT	M='L4'
XDOT59	G28_27	P28_27	G30_29	P30_29	G30_27	P30_27	DOT	M='L4'
XDOT60	G29_28	P29_28	G31_30	P31_30	G31_28	P31_28	DOT	M='L4'

*level 3 signal
XDOT61	G0	P0	G4_1	P4_1	G4_0	P4_0	DOT	M='L5'
XDOT62	G1_0	P1_0	G5_2	P5_2	G5_0	P5_0	DOT	M='L5'
XDOT63	G2_0	P2_0	G6_3	P6_3	G6_0	P6_0	DOT	M='L5'
XDOT64	G3_0	P3_0	G7_4	P7_4	G7_0	P7_0	DOT	M='L5'
XDOT65	G4_1	P4_1	G8_5	P8_5	G8_1	P8_1	DOT	M='L5'
XDOT66	G5_2	P5_2	G9_6	P9_6	G9_2	P9_2	DOT	M='L5'
XDOT67	G6_3	P6_3	G10_7	P10_7	G10_3	P10_3	DOT	M='L5'
XDOT68	G7_4	P7_4	G11_8	P11_8	G11_4	P11_4	DOT	M='L5'
XDOT69	G8_5	P8_5	G12_9	P12_9	G12_5	P12_5	DOT	M='L5'
XDOT70	G9_6	P9_6	G13_10	P13_10	G13_6	P13_6	DOT	M='L5'
XDOT71	G10_7	P10_7	G14_11	P14_11	G14_7	P14_7	DOT	M='L5'
XDOT72	G11_8	P11_8	G15_12	P15_12	G15_8	P15_8	DOT	M='L5'
XDOT73	G12_9	P12_9	G16_13	P16_13	G16_9	P16_9	DOT	M='L5'
XDOT74	G13_10	P13_10	G17_14	P17_14	G17_10	P17_10	DOT	M='L5'
XDOT75	G14_11	P14_11	G18_15	P18_15	G18_11	P18_11	DOT	M='L5'
XDOT76	G15_12	P15_12	G19_16	P19_16	G19_12	P19_12	DOT	M='L5'
XDOT77	G16_13	P16_13	G20_17	P20_17	G20_13	P20_13	DOT	M='L5'
XDOT78	G17_14	P17_14	G21_18	P21_18	G21_14	P21_14	DOT	M='L5'
XDOT79	G18_15	P18_15	G22_19	P22_19	G22_15	P22_15	DOT	M='L5'
XDOT80	G19_16	P19_16	G23_20	P23_20	G23_16	P23_16	DOT	M='L5'
XDOT81	G20_17	P20_17	G24_21	P24_21	G24_17	P24_17	DOT	M='L5'
XDOT82	G21_18	P21_18	G25_22	P25_22	G25_18	P25_18	DOT	M='L5'
XDOT83	G22_19	P22_19	G26_23	P26_23	G26_19	P26_19	DOT	M='L5'
XDOT84	G23_20	P23_20	G27_24	P27_24	G27_20	P27_20	DOT	M='L5'
XDOT85	G24_21	P24_21	G28_25	P28_25	G28_21	P28_21	DOT	M='L5'
XDOT86	G25_22	P25_22	G29_26	P29_26	G29_22	P29_22	DOT	M='L5'
XDOT87	G26_23	P26_23	G30_27	P30_27	G30_23	P30_23	DOT	M='L5'
XDOT88	G27_24	P27_24	G31_28	P31_28	G31_24	P31_24	DOT	M='L5'

*level 4 signal
XDOT89	G0	P0	G8_1	P8_1	G8_0	P8_0	DOT	M='L6'
XDOT90	G1_0	P1_0	G9_2	P9_2	G9_0	P9_0	DOT	M='L6'
XDOT91	G2_0	P2_0	G10_3	P10_3	G10_0	P10_0	DOT	M='L6'
XDOT92	G3_0	P3_0	G11_4	P11_4	G11_0	P11_0	DOT	M='L6'
XDOT93	G4_0	P4_0	G12_5	P12_5	G12_0	P12_0	DOT	M='L6'
XDOT94	G5_0	P5_0	G13_6	P13_6	G13_0	P13_0	DOT	M='L6'
XDOT95	G6_0	P6_0	G14_7	P14_7	G14_0	P14_0	DOT	M='L6'
XDOT96	G7_0	P7_0	G15_8	P15_8	G15_0	P15_0	DOT	M='L6'
XDOT97	G8_1	P8_1	G16_9	P16_9	G16_1	P16_1	DOT	M='L6'
XDOT98	G9_2	P9_2	G17_10	P17_10	G17_2	P17_2	DOT	M='L6'
XDOT99	G10_3	P10_3	G18_11	P18_11	G18_3	P18_3	DOT	M='L6'
XDOT100	G11_4	P11_4	G19_12	P19_12	G19_4	P19_4	DOT	M='L6'
XDOT101	G12_5	P12_5	G20_13	P20_13	G20_5	P20_5	DOT	M='L6'
XDOT102	G13_6	P13_6	G21_14	P21_14	G21_6	P21_6	DOT	M='L6'
XDOT103	G14_7	P14_7	G22_15	P22_15	G22_7	P22_7	DOT	M='L6'
XDOT104	G15_8	P15_8	G23_16	P23_16	G23_8	P23_8	DOT	M='L6'
XDOT105	G16_9	P16_9	G24_17	P24_17	G24_9	P24_9	DOT	M='L6'
XDOT106	G17_10	P17_10	G25_18	P25_18	G25_10	P25_10	DOT	M='L6'
XDOT107	G18_11	P18_11	G26_19	P26_19	G26_11	P26_11	DOT	M='L6'
XDOT108	G19_12	P19_12	G27_20	P27_20	G27_12	P27_12	DOT	M='L6'
XDOT109	G20_13	P20_13	G28_21	P28_21	G28_13	P28_13	DOT	M='L6'
XDOT110	G21_14	P21_14	G29_22	P29_22	G29_14	P29_14	DOT	M='L6'
XDOT111	G22_15	P22_15	G30_23	P30_23	G30_15	P30_15	DOT	M='L6'
XDOT112	G23_16	P23_16	G31_24	P31_24	G31_16	P31_16	DOT	M='L6'

*level 5 signal
XODT113	G0	P0	G16_1	P16_1	G16_0	P16_0	DOT	M='L7'
XDOT114	G1_0	P1_0	G17_2	P17_2	G17_0	P17_0	DOT	M='L7'
XDOT115	G2_0	P2_0	G18_3	P18_3	G18_0	P18_0	DOT	M='L7'
XDOT116	G3_0	P3_0	G19_4	P19_4	G19_0	P19_0	DOT	M='L7'
XDOT117	G4_0	P4_0	G20_5	P20_5	G20_0	P20_0	DOT	M='L7'
XDOT118	G5_0	P5_0	G21_6	P21_6	G21_0	P21_0	DOT	M='L7'
XDOT119	G6_0	P6_0	G22_7	P22_7	G22_0	P22_0	DOT	M='L7'
XDOT120	G7_0	P7_0	G23_8	P23_8	G23_0	P23_0	DOT	M='L7'
XDOT121	G8_0	P8_0	G24_9	P24_9	G24_0	P24_0	DOT	M='L7'
XDOT122	G9_0	P9_0	G25_10	P25_10	G25_0	P25_0	DOT	M='L7'
XDOT123	G10_0	P10_0	G26_11	P26_11	G26_0	P26_0	DOT	M='L7'
XDOT124	G11_0	P11_0	G27_12	P27_12	G27_0	P27_0	DOT	M='L7'
XDOT125	G12_0	P12_0	G28_13	P28_13	G28_0	P28_0	DOT	M='L7'
XDOT126	G13_0	P13_0	G29_14	P29_14	G29_0	P29_0	DOT	M='L7'
XDOT127	G14_0	P14_0	G30_15	P30_15	G30_0	P30_0	DOT	M='L7'
XDOT128	G15_0	P15_0	G31_16	P31_16	G31_0	P31_0	DOT	M='L7'

*sum genetation
XSUM0	A0	BO	S0	XOR2	M='L8'
XSUM1	P1	G0	S1	XOR2	M='L8'
XSUM2	P2	G1_0	S2	XOR2	M='L8'
XSUM3	P3	G2_0	S3	XOR2	M='L8'
XSUM4	P4	G3_0	S4	XOR2	M='L8'
XSUM5	P5	G4_0	S5	XOR2	M='L8'
XSUM6	P6	G5_0	S6	XOR2	M='L8'
XSUM7	P7	G6_0	S7	XOR2	M='L8'
XSUM8	P8	G7_0	S8	XOR2	M='L8'
XSUM9	P9	G8_0	S9	XOR2	M='L8'
XSUM10	P10	G9_0	S10	XOR2	M='L8'
XSUM11	P11	G10_0	S11	XOR2	M='L8'
XSUM12	P12	G11_0	S12	XOR2	M='L8'
XSUM13	P13	G12_0	S13	XOR2	M='L8'
XSUM14	P14	G13_0	S14	XOR2	M='L8'
XSUM15	P15	G14_0	S15	XOR2	M='L8'
XSUM16	P16	G15_0	S16	XOR2	M='L8'
XSUM17	P17	G16_0	S17	XOR2	M='L8'
XSUM18	P18	G17_0	S18	XOR2	M='L8'
XSUM19	P19	G18_0	S19	XOR2	M='L8'
XSUM20	P20	G19_0	S20	XOR2	M='L8'
XSUM21	P21	G20_0	S21	XOR2	M='L8'
XSUM22	P22	G21_0	S22	XOR2	M='L8'
XSUM23	P23	G22_0	S23	XOR2	M='L8'
XSUM24	P24	G23_0	S24	XOR2	M='L8'
XSUM25	P25	G24_0	S25	XOR2	M='L8'
XSUM26	P26	G25_0	S26	XOR2	M='L8'
XSUM27	P27	G26_0	S27	XOR2	M='L8'
XSUM28	P28	G27_0	S28	XOR2	M='L8'
XSUM29	P29	G28_0	S29	XOR2	M='L8'
XSUM30	P30	G29_0	S30	XOR2	M='L8'
XSUM31	P31	G30_0	S31	XOR2	M='L8'
.end
